`include "register_interface/typedef.svh"
`include "register_interface/assign.svh"

//typedef struct           packed {
//	 logic                 req;
//	 logic [31:0]          add;
//	 logic                 wen;
//	 logic [31:0]          wdata;
//	 logic [3:0]           be;
//} tcdm_req_t;
//typedef struct           packed {
//	 logic                 gnt;
//	 logic                 r_opc;
//	 logic [31:0]          r_rdata;
//	 logic                 r_valid;
//}tcdm_rsp_t;

module compute_output_wrapper
  import cutie_pkg::*;
  #(
    parameter int unsigned  TCDM_ADDR_WIDTH = 32,
    parameter int unsigned  TCDM_DATA_WIDTH = 32,
    parameter int unsigned TCDM_BE_WIDTH = TCDM_DATA_WIDTH/8,
    parameter int unsigned  TCDM_AUX_WIDTH = TCDM_DATA_WIDTH/8,

    parameter K = cutie_params::K,
    parameter N_I = cutie_params::N_I,
    parameter N_O = cutie_params::N_O,
    parameter IMAGEWIDTH = cutie_params::IMAGEWIDTH,
    parameter IMAGEHEIGHT = cutie_params::IMAGEHEIGHT,
    parameter WEIGHT_STAGGER = cutie_params::WEIGHT_STAGGER,
    parameter NUMACTMEMBANKSETS = cutie_params::NUMACTMEMBANKSETS,
    parameter WEIGHTBANKDEPTH = cutie_params::WEIGHTBANKDEPTH,
    parameter int unsigned  BANKSETSBITWIDTH = NUMACTMEMBANKSETS > 1 ? $clog2(NUMACTMEMBANKSETS) : 1,
    parameter int unsigned  NUMBANKS = K*WEIGHT_STAGGER,
    parameter int unsigned  TOTNUMTRITS = IMAGEWIDTH*IMAGEHEIGHT*N_I,
    parameter int unsigned  TRITSPERBANK = (TOTNUMTRITS+NUMBANKS-1)/NUMBANKS,
    parameter int unsigned  EFFECTIVETRITSPERWORD = N_I/WEIGHT_STAGGER,
    parameter int unsigned  PHYSICALTRITSPERWORD = ((EFFECTIVETRITSPERWORD + 4) / 5) * 5,
    parameter int unsigned  PHYSICALBITSPERWORD = PHYSICALTRITSPERWORD / 5 * 8,
    parameter int unsigned  ACTMEMBANKDEPTH = (TRITSPERBANK+EFFECTIVETRITSPERWORD-1)/EFFECTIVETRITSPERWORD,
    parameter int unsigned  ACTMEMFULLADDRESSBITWIDTH = $clog2(NUMBANKS*ACTMEMBANKDEPTH),
    parameter int unsigned  WEIGHTMEMFULLADDRESSBITWIDTH = $clog2(WEIGHTBANKDEPTH),
    parameter int unsigned  NUMENCODERS = PHYSICALBITSPERWORD/10
    )
   (
    input logic  soc_clk_i,
    input logic  soc_rst_ni,

    input logic  cutie_clk_i,
    input logic  cutie_rst_ni,

    input logic  cutie_memsleep_i,
    input logic  cutie_memgate_i,

    input logic  cutie_events_i,
    output logic cutie_events_o,

    input        tcdm_req_t tcdm_req_i,
    output       tcdm_rsp_t tcdm_rsp_o,
    input        reg_req_t reg_req_i,
    output       reg_rsp_t reg_rsp_o


    );

   import layer_params_reg_pkg::*;
   import cutie_params::*;

   //Convert the REG_BUS interface to the struct signals used by the autogenerated interface
   // typedef logic [31:0] data_t;
   // typedef logic [31:0] addr_t;
   // typedef logic [7:0]  strb_t;
   // `REG_BUS_TYPEDEF_REQ(reg_req_t, addr_t, data_t, strb_t)
   // `REG_BUS_TYPEDEF_RSP(reg_rsp_t, data_t)

   // Define REG_BUS interfaces on SoC clock domain side
   REG_BUS #(.ADDR_WIDTH(32), .DATA_WIDTH(32)) reg_bus(soc_clk_i);

   // each clock domain REG_BUS has a req channel and a rsp channel
   reg_req_t soc_domain_req, cutie_domain_req;
   reg_rsp_t soc_domain_rsp, cutie_domain_rsp;

   assign soc_domain_req = reg_req_i;
   assign reg_rsp_o = soc_domain_rsp;

   // // Convert APB to REB_BUS interface
   // apb_to_reg i_apb_to_reg
   //   (
   //    .clk_i(soc_clk_i),
   //    .rst_ni(soc_rst_ni),

   //    .penable_i(apb_penable_i),
   //    .pwrite_i(apb_pwrite_i),
   //    .paddr_i(apb_paddr_i),
   //    .psel_i(apb_psel_i),
   //    .pwdata_i(apb_pwdata_i),
   //    .prdata_o(apb_prdata_o),
   //    .pready_o(apb_pready_o),
   //    .pslverr_o(apb_pslverr_o),
   //    .reg_o(reg_bus)
   //    );

   // // REG_BUS interface to req and rsp channel structs
   // // This is done because the REG_CDC module only understands structs
   // `REG_BUS_ASSIGN_TO_REQ(soc_domain_req, reg_bus);
   // `REG_BUS_ASSIGN_FROM_RSP(reg_bus, soc_domain_rsp);

   reg_cdc #(.req_t(reg_req_t),.rsp_t(reg_rsp_t))
   i_reg_cdc(.src_clk_i(soc_clk_i),
	     .src_rst_ni(soc_rst_ni),
	     .src_req_i(soc_domain_req),
	     .src_rsp_o(soc_domain_rsp),
	     .dst_clk_i(cutie_clk_i),
	     .dst_rst_ni(cutie_rst_ni),
	     .dst_req_o(cutie_domain_req),
	     .dst_rsp_i(cutie_domain_rsp));

   layer_params_reg2hw_t reg_file_to_ip;
   layer_params_hw2reg_t ip_to_reg_file;

   layer_params_reg_top
     #(.reg_req_t(reg_req_t),
       .reg_rsp_t(reg_rsp_t))
   i_layer_params_reg_top
     (.clk_i(cutie_clk_i),
      .rst_ni(cutie_rst_ni),
      .reg_req_i(cutie_domain_req),
      .reg_rsp_o(cutie_domain_rsp),
      .reg2hw(reg_file_to_ip),
      .hw2reg(ip_to_reg_file),
      .devmode_i(1'b1)
      );

   logic                                    ctrl_valid_q;
   logic                                    threshold_qe_q;
   logic unsigned [$clog2(N_O):0]           layer_no_q;
   logic unsigned [$clog2(N_O):0]           layer_cnt_q, layer_cnt_d;
   logic [0:N_O-1]                          store_to_threshold;
   logic                                    thresh_fill_up_with_zeros_q, thresh_fill_up_with_zeros_d;
   logic                                    compute_done, compute_done_q;
   logic                                    start_compute_event;
   logic [0:N_O-1][$clog2(K*K*N_I):0]       fp_output;

   edge_propagator i_edge_prop_events_out
     (
      .clk_tx_i(cutie_clk_i),
      .rstn_tx_i(cutie_rst_ni),
      .edge_i(!compute_done_q && compute_done),
      .clk_rx_i(soc_clk_i),
      .rstn_rx_i(soc_rst_ni),
      .edge_o(cutie_events_o)
      );

   edge_propagator i_edge_prop_events_in
     (
      .clk_tx_i(soc_clk_i),
      .rstn_tx_i(soc_rst_ni),
      .edge_i(cutie_events_i),
      .clk_rx_i(cutie_clk_i),
      .rstn_rx_i(cutie_rst_ni),
      .edge_o(start_compute_event)
      );

   // assign ip_to_reg_file.fp_out = fp_output;

   always_comb begin

      if (start_compute_event) begin
	 ip_to_reg_file.ctrl2.d = 1'b0;
	 ip_to_reg_file.ctrl2.de = 1'b1;
      end else begin
	 ip_to_reg_file.ctrl2.d = 1'b0;
	 ip_to_reg_file.ctrl2.de = 1'b0;
      end

      for (int i = 0; i < N_O; i++) begin
	 ip_to_reg_file.fp_out[i] = fp_output[i];
      end

      store_to_threshold = '0;
      thresh_fill_up_with_zeros_d = 1'b0;

      layer_cnt_d = layer_cnt_q;

      if (reg_file_to_ip.ctrl1 && !ctrl_valid_q) begin
	 layer_cnt_d = 0;
      end

      ip_to_reg_file.thresholds.th_low.de = 1'b0;
      ip_to_reg_file.thresholds.th_low.d = '0;
      ip_to_reg_file.thresholds.th_high.de = 1'b0;
      ip_to_reg_file.thresholds.th_high.d = '0;

      if (!threshold_qe_q &&
	  reg_file_to_ip.thresholds.th_low.qe &&
	  reg_file_to_ip.thresholds.th_high.qe) begin
	 layer_cnt_d = layer_cnt_q + 1;
	 store_to_threshold = '0;
	 store_to_threshold[layer_cnt_q] = 1'b1;
      end else if (!reg_file_to_ip.ctrl1 && ctrl_valid_q) begin
	 ip_to_reg_file.thresholds.th_low.de = 1'b1;
	 ip_to_reg_file.thresholds.th_low.d = '0;
	 ip_to_reg_file.thresholds.th_high.de = 1'b1;
	 ip_to_reg_file.thresholds.th_high.d = '0;
	 thresh_fill_up_with_zeros_d = 1'b1;
      end

      if (thresh_fill_up_with_zeros_q) begin
	 store_to_threshold = {N_O{1'b1}} >> layer_cnt_q;
      end

      if(!compute_done_q && compute_done) begin
	 ip_to_reg_file.ctrl3.de = 1'b1;
	 ip_to_reg_file.ctrl3.d = 1'b1;
      end else begin
	 ip_to_reg_file.ctrl3.de = 1'b0;
	 ip_to_reg_file.ctrl3.d = 1'b0;
      end
   end

   always_ff @(posedge cutie_clk_i, negedge cutie_rst_ni) begin
      if(~cutie_rst_ni) begin
	 ctrl_valid_q <= 1'b0;
	 threshold_qe_q <= 1'b0;
	 layer_no_q <= '0;
	 layer_cnt_q <= '0;
	 compute_done_q <= '0;
	 thresh_fill_up_with_zeros_q <= '0;
      end else begin
	 ctrl_valid_q <= reg_file_to_ip.ctrl1;
	 threshold_qe_q <= (reg_file_to_ip.thresholds.th_low.qe &&
			    reg_file_to_ip.thresholds.th_high.qe);
	 layer_no_q <= reg_file_to_ip.feature_map.n_o;
	 layer_cnt_q <= layer_cnt_d;
	 compute_done_q <= compute_done;
	 thresh_fill_up_with_zeros_q <= thresh_fill_up_with_zeros_d;
      end
   end // always_ff @ (posedge clk_i, negedge rst_ni)

   logic [BANKSETSBITWIDTH-1:0]                actmem_bank_set;
   logic                                       actmem_we;
   logic                                       actmem_req;
   logic [ACTMEMFULLADDRESSBITWIDTH-1:0]       actmem_addr;
   logic [PHYSICALBITSPERWORD-1:0]             actmem_wdata;
   logic [PHYSICALBITSPERWORD-1:0]             actmem_rdata;
   logic                                       actmem_valid;
   logic [$clog2(N_O)-1:0]                     weightmem_bank;
   logic                                       weightmem_we;
   logic                                       weightmem_req;
   logic [WEIGHTMEMFULLADDRESSBITWIDTH-1:0]    weightmem_addr;
   logic [PHYSICALBITSPERWORD-1:0]             weightmem_wdata;
   logic [PHYSICALBITSPERWORD-1:0]             weightmem_rdata;
   logic                                       weightmem_valid;

   XBAR_TCDM_BUS cutie_tcdm_master();

   // TCDM Slave inputs
   assign cutie_tcdm_master.req = tcdm_req_i.req;
   assign cutie_tcdm_master.add = tcdm_req_i.add;
   assign cutie_tcdm_master.wen = tcdm_req_i.wen;
   assign cutie_tcdm_master.wdata = tcdm_req_i.wdata;
   assign cutie_tcdm_master.be = tcdm_req_i.be;

   // TCDM Slave outputs
   assign tcdm_rsp_o.gnt = cutie_tcdm_master.gnt;
   assign tcdm_rsp_o.r_valid = cutie_tcdm_master.r_valid;
   assign tcdm_rsp_o.r_rdata = cutie_tcdm_master.r_rdata;
   assign tcdm_rsp_o.r_opc = cutie_tcdm_master.r_opc;

   tcdm_to_mem i_tcdm_to_mem
   (/*AUTOINST*/
    // Interfaces
    .tcdm_slave                         (cutie_tcdm_master),
    // Outputs
    .actmem_bank_set_o                  (actmem_bank_set),
    .actmem_we_o                        (actmem_we),
    .actmem_req_o                       (actmem_req),
    .actmem_addr_o                      (actmem_addr),
    .actmem_wdata_o                     (actmem_wdata),
    .weightmem_bank_o                   (weightmem_bank),
    .weightmem_we_o                     (weightmem_we),
    .weightmem_req_o                    (weightmem_req),
    .weightmem_addr_o                   (weightmem_addr),
    .weightmem_wdata_o                  (weightmem_wdata),

    // Inputs
    .soc_clk_i                          (soc_clk_i),
    .soc_rst_ni                         (soc_rst_ni),
    .cutie_clk_i                        (cutie_clk_i),
    .cutie_rst_ni                       (cutie_rst_ni),
    .actmem_rdata_i                     (actmem_rdata),
    .actmem_valid_i                     (actmem_valid),
    .weightmem_rdata_i                  (weightmem_rdata),
    .weightmem_valid_i                  (weightmem_valid));


   cutie_top i_compute_output
     (// Outputs
      .actmem_external_acts_o(actmem_rdata),
      .actmem_external_valid_o(actmem_valid),
      .weightmem_external_weights_o(weightmem_rdata),
      .weightmem_external_valid_o(weightmem_valid),
      .compute_done_o     (compute_done),
      .fp_output_o(fp_output),
      // Inputs
      .clk_i              (cutie_clk_i),
      .rst_ni             (cutie_rst_ni),
      .actmem_external_bank_set_i(actmem_bank_set),
      .actmem_external_we_i(actmem_we),
      .actmem_external_req_i(actmem_req),
      .actmem_external_addr_i(actmem_addr),
      .actmem_external_wdata_i(actmem_wdata),
      .weightmem_external_bank_i(weightmem_bank),
      .weightmem_external_we_i(weightmem_we),
      .weightmem_external_req_i(weightmem_req),
      .weightmem_external_addr_i(weightmem_addr),
      .weightmem_external_wdata_i(weightmem_wdata),
      .ocu_thresh_pos_i   (reg_file_to_ip.thresholds.th_high.q),
      .ocu_thresh_neg_i   (reg_file_to_ip.thresholds.th_low.q),
      .ocu_thresholds_save_enable_i(store_to_threshold),
      .LUCA_store_to_fifo_i(!ctrl_valid_q && reg_file_to_ip.ctrl1),
      .LUCA_layer_imagewidth_i(reg_file_to_ip.feature_map.width),
      .LUCA_layer_imageheight_i(reg_file_to_ip.feature_map.height),
      .LUCA_layer_k_i     (reg_file_to_ip.kernel.k),
      .LUCA_layer_ni_i    (reg_file_to_ip.feature_map.n_i),
      .LUCA_layer_no_i    (reg_file_to_ip.feature_map.n_o),
      .LUCA_layer_stride_width_i(reg_file_to_ip.kernel.stride_w),
      .LUCA_layer_stride_height_i(reg_file_to_ip.kernel.stride_h),
      .LUCA_layer_padding_type_i(reg_file_to_ip.kernel.padding),
      .LUCA_pooling_enable_i(reg_file_to_ip.pooling.en),
      .LUCA_pooling_pooling_type_i(reg_file_to_ip.pooling.p_type),
      .LUCA_pooling_kernel_i(reg_file_to_ip.pooling.kernel),
      .LUCA_pooling_padding_type_i(reg_file_to_ip.pooling.padding),
      .LUCA_layer_skip_in_i('0),
      .LUCA_layer_skip_out_i('0),
      .LUCA_layer_is_tcn_i(reg_file_to_ip.tcn.is_tcn),
      .LUCA_layer_tcn_width_i(reg_file_to_ip.tcn.tcn_width),
      .LUCA_layer_tcn_width_mod_dil_i(reg_file_to_ip.tcn.tcn_width_mod_dil),
      .LUCA_layer_tcn_k_i (reg_file_to_ip.tcn.tcn_k),
      .LUCA_compute_disable_i(reg_file_to_ip.ctrl2)
      );

endmodule
